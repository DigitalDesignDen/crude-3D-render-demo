library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

PACKAGE vector_math_pkg IS
PROCEDURE SQ(SIGNAL Xcur, Ycur, Xpos, Ypos: IN INTEGER; SIGNAL RGB: OUT STD_LOGIC_VECTOR(9 downto 0); SIGNAL DRAW: OUT STD_LOGIC);
PROCEDURE DIFF(VARIABLE X1, Y1, X2, Y2: IN INTEGER; VARIABLE dX,dY: OUT INTEGER);
PROCEDURE DET(VARIABLE X1,Y1,X2,Y2: IN INTEGER; VARIABLE LINEAR_DEPENDENT: OUT BOOLEAN);
END vector_math_pkg;

PACKAGE BODY vector_math_pkg IS
PROCEDURE SQ(SIGNAL Xcur, Ycur, Xpos, Ypos: IN INTEGER; SIGNAL RGB: OUT STD_LOGIC_VECTOR(9 downto 0); SIGNAL DRAW: OUT STD_LOGIC) IS
BEGIN

IF Xcur>Xpos AND Xcur<(Xpos+100) AND Ycur>Ypos AND Ycur<(Ypos+100) THEN
	RGB <= "0000000111";
	DRAW <= '1';
ELSE
	DRAW <= '0';
END IF;

END SQ;

PROCEDURE DIFF(X1, Y1, X2, Y2: IN INTEGER; dX,dY: OUT INTEGER) IS
BEGIN
dX :=  X1 - X2;
dY :=  Y1 - Y2;
END DIFF;

PROCEDURE DET(X1,Y1,X2,Y2 : IN INTEGER; LINEAR_DEPENDENT : OUT BOOLEAN) IS
BEGIN

IF((X1 * Y2) - (Y1 * X2) >= -30 AND (X1 * Y2) - (Y1 * X2) <= 30) THEN
	LINEAR_DEPENDENT :=  TRUE;
ELSE
	LINEAR_DEPENDENT :=  FALSE;
END IF;
END DET;
END vector_math_pkg;